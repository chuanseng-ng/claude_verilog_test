// rv32i_decode.sv
// RV32I Instruction Decoder

module rv32i_decode (
  // Instruction input
  input  logic [31:0] instruction,

  // Decoded register addresses
  output logic [4:0]  rs1,        // Source register 1
  output logic [4:0]  rs2,        // Source register 2
  output logic [4:0]  rd,         // Destination register

  // ALU control
  output logic [3:0]  alu_op,     // ALU operation (using approved encoding)
  output logic [1:0]  alu_src_a,  // ALU operand A select: 00=rs1, 01=PC, 10=zero
  output logic        alu_src_b,  // 0=rs2, 1=immediate

  // Immediate format
  output logic [2:0]  imm_fmt,    // Immediate format for imm_gen

  // Register file control
  output logic        reg_wr_en,  // Register write enable

  // Memory control
  output logic        mem_rd,     // Memory read enable
  output logic        mem_wr,     // Memory write enable
  output logic [2:0]  mem_size,   // 000=byte, 001=half, 010=word
  output logic        mem_unsigned, // Unsigned load

  // Branch/Jump control
  output logic        branch,     // Branch instruction
  output logic [2:0]  branch_op,  // Branch comparison type
  output logic        jump,       // Jump instruction (JAL/JALR)
  output logic        jalr,       // JALR (PC-relative vs register-relative)

  // Control signals
  output logic        pc_src,     // 0=PC+4, 1=branch/jump target
  output logic        illegal,    // Illegal instruction flag
  output logic        ebreak      // EBREAK instruction (triggers CPU halt)
);

  // Extract instruction fields
  logic [6:0] opcode;
  logic [2:0] funct3;
  logic [6:0] funct7;

  assign opcode = instruction[6:0];
  assign funct3 = instruction[14:12];
  assign funct7 = instruction[31:25];
  assign rs1    = instruction[19:15];
  assign rs2    = instruction[24:20];
  assign rd     = instruction[11:7];

  // Opcode definitions (RV32I)
  localparam [6:0] OP_LUI    = 7'b0110111;
  localparam [6:0] OP_AUIPC  = 7'b0010111;
  localparam [6:0] OP_JAL    = 7'b1101111;
  localparam [6:0] OP_JALR   = 7'b1100111;
  localparam [6:0] OP_BRANCH = 7'b1100011;
  localparam [6:0] OP_LOAD   = 7'b0000011;
  localparam [6:0] OP_STORE  = 7'b0100011;
  localparam [6:0] OP_IMM    = 7'b0010011;  // ALU immediate operations
  localparam [6:0] OP_REG    = 7'b0110011;  // ALU register operations
  localparam [6:0] OP_SYSTEM = 7'b1110011;  // SYSTEM instructions (EBREAK, ECALL)

  // Funct3 definitions for branches
  localparam [2:0] FUNCT3_BEQ  = 3'b000;
  localparam [2:0] FUNCT3_BNE  = 3'b001;
  localparam [2:0] FUNCT3_BLT  = 3'b100;
  localparam [2:0] FUNCT3_BGE  = 3'b101;
  localparam [2:0] FUNCT3_BLTU = 3'b110;
  localparam [2:0] FUNCT3_BGEU = 3'b111;

  // Funct3 definitions for loads
  localparam [2:0] FUNCT3_LB  = 3'b000;
  localparam [2:0] FUNCT3_LH  = 3'b001;
  localparam [2:0] FUNCT3_LW  = 3'b010;
  localparam [2:0] FUNCT3_LBU = 3'b100;
  localparam [2:0] FUNCT3_LHU = 3'b101;

  // Funct3 definitions for stores
  localparam [2:0] FUNCT3_SB = 3'b000;
  localparam [2:0] FUNCT3_SH = 3'b001;
  localparam [2:0] FUNCT3_SW = 3'b010;

  // Funct3 definitions for ALU operations
  localparam [2:0] FUNCT3_ADD_SUB = 3'b000;
  localparam [2:0] FUNCT3_SLL     = 3'b001;
  localparam [2:0] FUNCT3_SLT     = 3'b010;
  localparam [2:0] FUNCT3_SLTU    = 3'b011;
  localparam [2:0] FUNCT3_XOR     = 3'b100;
  localparam [2:0] FUNCT3_SRL_SRA = 3'b101;
  localparam [2:0] FUNCT3_OR      = 3'b110;
  localparam [2:0] FUNCT3_AND     = 3'b111;

  // ALU operation encodings (from approved scheme)
  localparam [3:0] ALU_ADD  = 4'b0000;
  localparam [3:0] ALU_SUB  = 4'b0001;
  localparam [3:0] ALU_SLL  = 4'b0010;
  localparam [3:0] ALU_SLT  = 4'b0011;
  localparam [3:0] ALU_SLTU = 4'b0100;
  localparam [3:0] ALU_XOR  = 4'b0101;
  localparam [3:0] ALU_SRL  = 4'b0110;
  localparam [3:0] ALU_SRA  = 4'b0111;
  localparam [3:0] ALU_OR   = 4'b1000;
  localparam [3:0] ALU_AND  = 4'b1001;

  // Immediate format encodings
  localparam [2:0] FMT_I = 3'b000;
  localparam [2:0] FMT_S = 3'b001;
  localparam [2:0] FMT_B = 3'b010;
  localparam [2:0] FMT_U = 3'b011;
  localparam [2:0] FMT_J = 3'b100;
  localparam [2:0] FMT_R = 3'b101;

  // ALU operand A source select encodings
  localparam [1:0] SRC_A_RS1  = 2'b00;  // Select rs1_data
  localparam [1:0] SRC_A_PC   = 2'b01;  // Select PC (for AUIPC)
  localparam [1:0] SRC_A_ZERO = 2'b10;  // Select zero (for LUI)

  // Main decoder logic
  always_comb begin
    // Default values (prevents latches)
    alu_op       = ALU_ADD;
    alu_src_a    = SRC_A_RS1;  // Default: rs1_data
    alu_src_b    = 1'b0;       // Default: rs2
    imm_fmt      = FMT_I;
    reg_wr_en    = 1'b0;
    mem_rd       = 1'b0;
    mem_wr       = 1'b0;
    mem_size     = 3'b010;  // Word
    mem_unsigned = 1'b0;
    branch       = 1'b0;
    branch_op    = 3'b000;
    jump         = 1'b0;
    jalr         = 1'b0;
    pc_src       = 1'b0;
    illegal      = 1'b0;
    ebreak       = 1'b0;

    case (opcode)
      // ================================================================
      // LUI - Load Upper Immediate
      // rd = imm[31:12] << 12 = 0 + U-immediate
      // ================================================================
      OP_LUI: begin
        imm_fmt   = FMT_U;
        reg_wr_en = 1'b1;
        alu_op    = ALU_ADD;
        alu_src_a = SRC_A_ZERO;  // Select zero operand
        alu_src_b = 1'b1;        // Select U-immediate
      end

      // ================================================================
      // AUIPC - Add Upper Immediate to PC
      // rd = PC + (imm[31:12] << 12)
      // ================================================================
      OP_AUIPC: begin
        imm_fmt   = FMT_U;
        reg_wr_en = 1'b1;
        alu_op    = ALU_ADD;
        alu_src_a = SRC_A_PC;  // Select PC
        alu_src_b = 1'b1;      // Select U-immediate
      end

      // ================================================================
      // JAL - Jump and Link
      // rd = PC + 4, PC = PC + imm
      // ================================================================
      OP_JAL: begin
        imm_fmt   = FMT_J;
        reg_wr_en = 1'b1;
        jump      = 1'b1;
        jalr      = 1'b0;
        // Need to save PC+4 to rd and update PC to PC+imm
      end

      // ================================================================
      // JALR - Jump and Link Register
      // rd = PC + 4, PC = (rs1 + imm) & ~1
      // ================================================================
      OP_JALR: begin
        if (funct3 == 3'b000) begin
          imm_fmt   = FMT_I;
          reg_wr_en = 1'b1;
          jump      = 1'b1;
          jalr      = 1'b1;
        end else begin
          illegal = 1'b1;  // Invalid funct3 for JALR
        end
      end

      // ================================================================
      // BRANCH - Conditional branches
      // BEQ, BNE, BLT, BGE, BLTU, BGEU
      // ================================================================
      OP_BRANCH: begin
        imm_fmt   = FMT_B;
        branch    = 1'b1;
        branch_op = funct3;

        case (funct3)
          FUNCT3_BEQ,
          FUNCT3_BNE,
          FUNCT3_BLT,
          FUNCT3_BGE,
          FUNCT3_BLTU,
          FUNCT3_BGEU: begin
            illegal = 1'b0;
          end
          default: begin
            illegal = 1'b1;  // Invalid branch type
          end
        endcase
      end

      // ================================================================
      // LOAD - Load instructions
      // LB, LH, LW, LBU, LHU
      // ================================================================
      OP_LOAD: begin
        imm_fmt   = FMT_I;
        reg_wr_en = 1'b1;
        mem_rd    = 1'b1;
        alu_op    = ALU_ADD;
        alu_src_a = 1'b0;  // rs1
        alu_src_b = 1'b1;  // Immediate

        case (funct3)
          FUNCT3_LB: begin
            mem_size     = 3'b000;  // Byte
            mem_unsigned = 1'b0;    // Signed
          end
          FUNCT3_LH: begin
            mem_size     = 3'b001;  // Halfword
            mem_unsigned = 1'b0;    // Signed
          end
          FUNCT3_LW: begin
            mem_size     = 3'b010;  // Word
            mem_unsigned = 1'b0;    // Don't care for word
          end
          FUNCT3_LBU: begin
            mem_size     = 3'b000;  // Byte
            mem_unsigned = 1'b1;    // Unsigned
          end
          FUNCT3_LHU: begin
            mem_size     = 3'b001;  // Halfword
            mem_unsigned = 1'b1;    // Unsigned
          end
          default: begin
            illegal = 1'b1;
          end
        endcase
      end

      // ================================================================
      // STORE - Store instructions
      // SB, SH, SW
      // ================================================================
      OP_STORE: begin
        imm_fmt   = FMT_S;
        mem_wr    = 1'b1;
        alu_op    = ALU_ADD;
        alu_src_a = 1'b0;  // rs1
        alu_src_b = 1'b1;  // Immediate

        case (funct3)
          FUNCT3_SB: begin
            mem_size = 3'b000;  // Byte
          end
          FUNCT3_SH: begin
            mem_size = 3'b001;  // Halfword
          end
          FUNCT3_SW: begin
            mem_size = 3'b010;  // Word
          end
          default: begin
            illegal = 1'b1;
          end
        endcase
      end

      // ================================================================
      // OP_IMM - Immediate ALU operations
      // ADDI, SLTI, SLTIU, XORI, ORI, ANDI, SLLI, SRLI, SRAI
      // ================================================================
      OP_IMM: begin
        imm_fmt   = FMT_I;
        reg_wr_en = 1'b1;
        alu_src_a = 1'b0;  // rs1
        alu_src_b = 1'b1;  // Immediate

        case (funct3)
          FUNCT3_ADD_SUB: begin
            alu_op = ALU_ADD;  // ADDI
          end
          FUNCT3_SLT: begin
            alu_op = ALU_SLT;  // SLTI
          end
          FUNCT3_SLTU: begin
            alu_op = ALU_SLTU;  // SLTIU
          end
          FUNCT3_XOR: begin
            alu_op = ALU_XOR;  // XORI
          end
          FUNCT3_OR: begin
            alu_op = ALU_OR;  // ORI
          end
          FUNCT3_AND: begin
            alu_op = ALU_AND;  // ANDI
          end
          FUNCT3_SLL: begin
            // SLLI - Check funct7 for validity
            if (funct7 == 7'b0000000) begin
              alu_op = ALU_SLL;
            end else begin
              illegal = 1'b1;
            end
          end
          FUNCT3_SRL_SRA: begin
            // SRLI or SRAI - distinguished by funct7[5]
            if (funct7 == 7'b0000000) begin
              alu_op = ALU_SRL;  // SRLI
            end else if (funct7 == 7'b0100000) begin
              alu_op = ALU_SRA;  // SRAI
            end else begin
              illegal = 1'b1;
            end
          end
          default: begin
            illegal = 1'b1;
          end
        endcase
      end

      // ================================================================
      // OP_REG - Register-register ALU operations
      // ADD, SUB, SLL, SLT, SLTU, XOR, SRL, SRA, OR, AND
      // ================================================================
      OP_REG: begin
        imm_fmt   = FMT_R;
        reg_wr_en = 1'b1;
        alu_src_a = 1'b0;  // rs1
        alu_src_b = 1'b0;  // rs2

        case (funct3)
          FUNCT3_ADD_SUB: begin
            // ADD or SUB - distinguished by funct7[5]
            if (funct7 == 7'b0000000) begin
              alu_op = ALU_ADD;  // ADD
            end else if (funct7 == 7'b0100000) begin
              alu_op = ALU_SUB;  // SUB
            end else begin
              illegal = 1'b1;
            end
          end
          FUNCT3_SLL: begin
            if (funct7 == 7'b0000000) begin
              alu_op = ALU_SLL;  // SLL
            end else begin
              illegal = 1'b1;
            end
          end
          FUNCT3_SLT: begin
            if (funct7 == 7'b0000000) begin
              alu_op = ALU_SLT;  // SLT
            end else begin
              illegal = 1'b1;
            end
          end
          FUNCT3_SLTU: begin
            if (funct7 == 7'b0000000) begin
              alu_op = ALU_SLTU;  // SLTU
            end else begin
              illegal = 1'b1;
            end
          end
          FUNCT3_XOR: begin
            if (funct7 == 7'b0000000) begin
              alu_op = ALU_XOR;  // XOR
            end else begin
              illegal = 1'b1;
            end
          end
          FUNCT3_SRL_SRA: begin
            // SRL or SRA - distinguished by funct7[5]
            if (funct7 == 7'b0000000) begin
              alu_op = ALU_SRL;  // SRL
            end else if (funct7 == 7'b0100000) begin
              alu_op = ALU_SRA;  // SRA
            end else begin
              illegal = 1'b1;
            end
          end
          FUNCT3_OR: begin
            if (funct7 == 7'b0000000) begin
              alu_op = ALU_OR;  // OR
            end else begin
              illegal = 1'b1;
            end
          end
          FUNCT3_AND: begin
            if (funct7 == 7'b0000000) begin
              alu_op = ALU_AND;  // AND
            end else begin
              illegal = 1'b1;
            end
          end
          default: begin
            illegal = 1'b1;
          end
        endcase
      end

      // ================================================================
      // SYSTEM - EBREAK instruction
      // EBREAK: opcode=0b1110011, funct3=0, imm12=1
      // Encoding: 0x00100073
      // ================================================================
      OP_SYSTEM: begin
        if (funct3 == 3'b000 && instruction[31:20] == 12'h001) begin
          // EBREAK - trigger CPU halt via debug interface
          ebreak    = 1'b1;
          illegal   = 1'b0;
          // No register write, no memory access
        end else begin
          // Other SYSTEM instructions (ECALL, CSR ops) not supported in Phase 1
          illegal = 1'b1;
        end
      end

      // ================================================================
      // Default - Illegal instruction
      // ================================================================
      default: begin
        illegal = 1'b1;
      end
    endcase
  end

endmodule

// ============================================================================
// HUMAN REVIEW CHECKLIST
// ============================================================================
//
// Please verify the following before approving this decoder:
//
// ✓ All 37 RV32I instructions are covered:
//   - Arithmetic: ADD, SUB, ADDI (3)
//   - Logical: AND, OR, XOR, ANDI, ORI, XORI (6)
//   - Shifts: SLL, SRL, SRA, SLLI, SRLI, SRAI (6)
//   - Compare: SLT, SLTU, SLTI, SLTIU (4)
//   - Branches: BEQ, BNE, BLT, BGE, BLTU, BGEU (6)
//   - Jumps: JAL, JALR (2)
//   - Loads: LB, LH, LW, LBU, LHU (5)
//   - Stores: SB, SH, SW (3)
//   - Upper: LUI, AUIPC (2)
//   TOTAL: 37 instructions
//
// ✓ Similar instructions properly distinguished:
//   - ADD vs SUB (funct7[5])
//   - SRL vs SRA (funct7[5])
//   - SRLI vs SRAI (funct7[5])
//   - LB vs LBU (funct3)
//   - LH vs LHU (funct3)
//
// ✓ Control signal encoding is correct and complete
//
// ✓ Illegal instruction detection covers:
//   - Invalid opcodes
//   - Invalid funct3/funct7 combinations
//   - Reserved encodings
//
// ✓ ALU operation encodings match approved scheme
//
// ✓ Immediate formats match RV32I specification
//
// ============================================================================
